//defining NOT gate
module v7404(pin1, pin3, pin5, pin9, pin11, pin13, pin2, pin4, pin6, pin8, pin10, pin12);

    input pin1, pin3, pin5, pin9, pin11, pin13;
    output pin2, pin4, pin6, pin8, pin10, pin12;

    assign pin2 = ~pin1;
    assign pin4 = ~pin3;
    assign pin6 = ~pin5;
    assign pin8 = ~pin9;
    assign pin10 = ~pin11;
    assign pin12 = ~pin13;
endmodule

//defining AND gate
module v7408(pin1, pin2, pin4, pin5, pin9, pin10, pin12, pin13, pin3, pin6, pin8, pin11);
   
    input pin1, pin2, pin4, pin5, pin9, pin10, pin12, pin13;
    output pin3, pin6, pin8, pin11;

    assign pin3 = pin1&pin2;
    assign pin6 = pin4&pin5;
    assign pin8 = pin9&pin10;
    assign pin11 = pin12&pin13;
endmodule

//defining OR gate
module v7432(pin1, pin2, pin4, pin5, pin9, pin10, pin12, pin13, pin3, pin6, pin8, pin11);

    input pin1, pin2, pin4, pin5, pin9, pin10, pin12, pin13;
    output pin3, pin6, pin8, pin11;

    assign pin3 = pin1|pin2;
    assign pin6 = pin4|pin5;
    assign pin8 = pin9|pin10;
    assign pin11 = pin12|pin13;
endmodule

//defining mux2to1
module mux2to1 (x,y,s,m);
    input x,y,s;
    output m;

    wire Connection1, Connection2, Connection3;

    v7404 notGate(
        .pin1(s), .pin2(Connection1)
    );

    v7408 andGate(
        .pin1(Connection1),
        .pin2(x),
        .pin3(Connection2),
        .pin4(s),
        .pin5(y),
        .pin6(Connection3)
    );

    v7432 orGate(
        .pin1(Connection2), .pin2(Connection3), .pin3(m)
    );

endmodule